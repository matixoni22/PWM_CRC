
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all


entity CRC-16_coder is
    Port ( In_coder : in  STD_LOGIC;
           Out_coder : out  STD_LOGIC;
           Out_crc : out  STD_LOGIC);
end CRC-16_coder;

architecture a_CRC-16 of CRC-16_coder is

begin


end a_CRC-16;

